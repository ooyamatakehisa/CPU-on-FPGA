module flopenableEX #(parameter WIDTH=8)
				(	
					input clk, reset,flush,
					input [WIDTH-1:0] d,
					output reg [WIDTH-1:0] q );
					
	always @ (posedge clk, posedge reset) begin
		if (reset) q <= 0;
		else if(flush) q <= 0 ;
		else 
			q <= d;
		end
	
endmodule